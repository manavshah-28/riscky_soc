import riscky_pkg::*;

module extender(
);

endmodule