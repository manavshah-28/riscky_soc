module instr_mem(
    input logic rst,
    input logic [],

);

endmodule