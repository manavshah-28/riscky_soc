package riscky_pkg;
parameter int XLEN = 64;
endpackage