import riscky_pkg::*;

module fetch(
    input clk, rst_n, PC_sel,
    input [XLEN-1:0] PC_target,
    output [ILEN-1:0] Instr

);

endmodule